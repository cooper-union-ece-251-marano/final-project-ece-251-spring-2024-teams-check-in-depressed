//////////////////////////////////////////////////////////////////////////////////
// The Cooper Union
// ECE 251 Spring 2024
// Engineer: Tiffany Shum & Lani Wang
// 
//     Create Date: 2024-05-08
//     Module Name: tb_alu
//     Description: Test bench for 16 bit ALU
//
// Revision: 1.0
//
//////////////////////////////////////////////////////////////////////////////////
`ifndef TB_ALU
`define TB_ALU

`timescale 1ns/100ps
`include "alu.sv"

module tb_alu;
    parameter n = 16;
    logic [(n-1):0] i1, i2;
    logic [2:0] op;
    logic zero;

    initial begin
		$dumpfile("alu.vcd");
        $dumpvars(0, uut);
      $monitor("i1 = %b i2 = %b opcode = %b", i1, i2, op);
    end

    initial begin
	    i1 <= 16'b0000000000000000;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b000;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;
        
	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b001;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b010;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b011;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b100;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b101;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b110;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;

	    #10 i1 <= 16'b0001000101000101;
	    i2 <= 16'b0000000000000000;
	    op <= 3'b111;
	    #10 i1 <= 16'b1111111111111111;
	    i2 <= 16'b1011011101111110;
	    #10 i1 <= 16'b0001000101000101;
	    #10 i1 <= 16'b0000000000000000;
    end

    alu uut(.i1(i1), .i2(i2), .op(op));

endmodule
`endif // TB_ALU